/**/
`include "C:/Users/hp/Desktop/my_1942/define.v"
module noiseWave (
    input byte0
);
    
endmodule