/*
    nameTableRam:名称表32x30的尺寸，一共960个title
*/

`include "C:/Users/hp/Desktop/my1942Game/RTL/src/game/PPU/define.v"
module nameTableRam(
    //cortex-m0
    input clk,
    input [`NAMETABLE_AHBBUS_ADDRWIDTH-1:0] addra,
    input [`NAMETABLE_AHBBUS_ADDRWIDTH-1:0] addrb,
    input [31:0] dina,
    input [3:0] wea,
    output reg [31:0] doutb,

    //到tiledraw函数
    input clk_tileDraw,
    input [`NAMETABLE_AHBBUS_ADDRWIDTH-1:0] nameTableRamIndex,
    output reg [31:0] nameTableRamDataO,
    input wire    [9-1:0]  attributeAddr, //0~32*30/4=240
    output reg    [4*(`BYTE)-1:0]     attributeTableDataO
);

    // (* ram_style="block" *) reg  [4*(`BYTE)-1:0] nameTableRam [0:((`NAMETABLE_HEIGHT)*(`NAMETABLE_WIDTH))>>2-1];
    (* ram_style="block" *) reg  [4*(`BYTE)-1:0] nameTableRam [0:512-1];//适配安路的板子进行的修改，与地址线的位宽保持一致
    initial begin
	    $readmemh("C:/Users/hp/Desktop/my1942Game/RTL/src/game/PPU/backGround/nameTable_test02.txt", nameTableRam);
	end

/*与CPU M0软核的交互 注意与其他的ram写的高低位位置不一样*/
    always@(posedge clk) begin
        if(wea[3]) nameTableRam[addra][7:0] <= dina[07:00];
    end
    always@(posedge clk) begin
        if(wea[2]) nameTableRam[addra][15:8] <= dina[15:08];
    end
    always@(posedge clk) begin
        if(wea[1]) nameTableRam[addra][23:16] <= dina[23:16];
    end
    always@(posedge clk) begin
        if(wea[0]) nameTableRam[addra][31:24] <= dina[31:24];
    end

    always@(posedge clk) begin
        doutb <= nameTableRam[addrb];
    end

/*与其他PPU模块的交互*/
    always@(posedge clk_tileDraw) begin
        nameTableRamDataO <= nameTableRam[nameTableRamIndex];
    end

    always@(posedge clk_tileDraw)begin
        attributeTableDataO<=nameTableRam[attributeAddr];
    end

endmodule